module encorder( out, in ) ;
  input [3:0] in ; 
  output [6:0] out ;

  assign out[6:0] = ( in[3:0] == 0 ) ? 7'b0111111 :
                    ( in[3:0] == 1 ) ? 7'b0000110 :
                    ( in[3:0] == 2 ) ? 7'b1011011 :
                    ( in[3:0] == 3 ) ? 7'b1001111 :
                    ( in[3:0] == 4 ) ? 7'b1100110 :
                    ( in[3:0] == 5 ) ? 7'b1101101 :
                    ( in[3:0] == 6 ) ? 7'b1111101 :
                    ( in[3:0] == 7 ) ? 7'b0100111 :
                    ( in[3:0] == 8 ) ? 7'b1111111 :
                    ( in[3:0] == 9 ) ? 7'b1101111 : 
                    ( in[3:0] == 10) ? 7'b1110111 : 
                    ( in[3:0] == 11) ? 7'b1111100 :
                    ( in[3:0] == 12) ? 7'b0111001 : 
                    ( in[3:0] == 13) ? 7'b1011110 :
                    ( in[3:0] == 14) ? 7'b1111001 :
                    ( in[3:0] == 15) ? 7'b1110001 : 7'b0000000 ;
                    
endmodule




