module cpu15(CLK, RESET_N, IO65_IN, IO65_OUT);
input           CLK;
input           RESET_N;
input   [15:0]  IO65_IN;
output  [15:0]  IO65_OUT;

// statement

endmodule